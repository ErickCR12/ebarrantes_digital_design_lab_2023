module videoGen(input logic [9:0] x, y,
					 output logic [7:0] r, g, b);

endmodule