module victory_tb();

	reg [6:0] tab [7:0][7:0];
	reg [7:0]bombas;
	logic clk, rst;
	
	
endmodule