library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

entity FullAdder4Bit_tb is -- no inputs or outputs
end FullAdder4Bit_tb;

architecture fulladder4bit_tb of FullAdder4Bit_tb is
	component FullAdder_4bit
		Port ( A : in STD_LOGIC_VECTOR(3 downto 0);
				 B : in STD_LOGIC_VECTOR(3 downto 0);
				 Cin : in STD_LOGIC;
				 Sum : out STD_LOGIC_VECTOR(3 downto 0);
				 Cout : out STD_LOGIC);
	end component;
	signal A, B : STD_LOGIC_VECTOR(3 downto 0);
	signal Cin : STD_LOGIC;
	signal Sum : STD_LOGIC_VECTOR(3 downto 0);
	signal Cout : STD_LOGIC;

begin
	-- Instancia del sumador
	UUT: FullAdder_4bit port map (A, B, Cin, Sum, Cout);
	process begin
		-- Establecer valores iniciales
		A <= "0000";
		B <= "0000";
		Cin <= '0';
		wait for 0.2 ns;

		-- Prueba 1
		A <= "0101";
		B <= "0010";
		Cin <= '0';
		wait for 0.2 ns;

		-- Prueba 2
		A <= "1100";
		B <= "1011";
		Cin <= '1';
		wait for 0.2 ns;

		-- Prueba 3
		A <= "1111";
		B <= "0001";
		Cin <= '0';
		wait for 0.2 ns;

		-- Prueba 4
		A <= "1010";
		B <= "0101";
		Cin <= '1';
		wait for 0.2 ns;

		-- Detener la simulación
		wait;
	end process;
end;