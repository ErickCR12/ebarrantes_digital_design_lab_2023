module decoBCD(A,B,C,D,a,b,c,d,e,f,g,h)

			input A,B,C,D
			output a,b,c,d,e,f,g,h
						always @(A,B,C,D)
				begin
				if(A==1'b0 & B==1'b0 & C==1'b0 & D==1'b0) a==1'b0

endmodule